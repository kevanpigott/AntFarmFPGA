//Author: Kevan Pigott
module only2quadrants(in,out);
input[1:0]in;
output [1:0]out =in[1];
endmodule