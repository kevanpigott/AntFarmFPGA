//Author:Kevan Pigott
module kevansVGAtesterthing(out);
output [104:0] out=131'hfffffffffffffffffffdfffffffffffff;





endmodule