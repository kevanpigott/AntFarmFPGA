//Author: Kevan Pigott
module errorSpacePush(outERROR);

output [11:0]outERROR=11'hff;

endmodule