//Author: Kevan Pigott
module quadrantDraw (outA,outB,outC,outD,outE);

output [0:20]outA=21'o1111717;
output [0:20]outB=21'o7771177;
output [0:20]outC=21'o7171717;
output [0:20]outD=21'o7771111;
output [0:20]outE=21'o1171111;

endmodule